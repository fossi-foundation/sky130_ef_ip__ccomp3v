magic
tech sky130A
magscale 1 2
timestamp 1747682096
<< dnwell >>
rect -127 6072 10341 10125
rect -127 -2512 11133 6072
<< nwell >>
rect -236 10017 10450 10234
rect -236 5932 79 10017
rect 10145 6344 10450 10017
rect 10246 6187 10450 6344
rect 5141 6186 10450 6187
rect -236 1870 101 5932
rect 5141 5929 11242 6186
rect 9361 5860 11242 5929
rect 10907 1870 11242 5860
rect -236 -2306 79 1870
rect 10927 -2306 11242 1870
rect -236 -2621 11242 -2306
<< mvpsubdiff >>
rect -358 10323 -298 10357
rect 10517 10323 10577 10357
rect -358 10297 -324 10323
rect 10543 10297 10577 10323
rect 10543 6313 10577 6344
rect 10543 6279 10615 6313
rect 11230 6279 11369 6313
rect 11335 6248 11369 6279
rect -358 -2712 -324 -2686
rect 11335 -2712 11369 -2686
rect -358 -2746 -298 -2712
rect 11309 -2746 11369 -2712
<< mvnsubdiff >>
rect -170 10148 10384 10168
rect -170 10114 -90 10148
rect 10304 10114 10384 10148
rect -170 10094 10384 10114
rect -170 10088 -96 10094
rect -170 -2475 -150 10088
rect -116 -2475 -96 10088
rect 10310 10088 10384 10094
rect 10310 6152 10330 10088
rect 10364 6152 10384 10088
rect 10310 6120 10384 6152
rect 10310 6101 11176 6120
rect 10310 6067 10364 6101
rect 11086 6072 11176 6101
rect 11086 6067 11122 6072
rect 10310 6046 11122 6067
rect -170 -2481 -96 -2475
rect 11102 -2466 11122 6046
rect 11156 -2466 11176 6072
rect 11102 -2481 11176 -2466
rect -170 -2501 11176 -2481
rect -170 -2535 -90 -2501
rect 11086 -2535 11176 -2501
rect -170 -2555 11176 -2535
<< mvpsubdiffcont >>
rect -298 10323 10517 10357
rect -358 -2686 -324 10297
rect 10543 6344 10577 10297
rect 10615 6279 11230 6313
rect 11335 -2686 11369 6248
rect -298 -2746 11309 -2712
<< mvnsubdiffcont >>
rect -90 10114 10304 10148
rect -150 -2475 -116 10088
rect 10330 6152 10364 10088
rect 10364 6067 11086 6101
rect 11122 -2466 11156 6072
rect -90 -2535 11086 -2501
<< locali >>
rect -358 10323 -298 10357
rect 10517 10323 10577 10357
rect -358 10317 10577 10323
rect -358 10297 -216 10317
rect -324 10268 -216 10297
rect 10415 10297 10577 10317
rect 10415 10268 10543 10297
rect -324 10235 10543 10268
rect -324 10154 -237 10235
rect -324 -2546 -312 10154
rect -260 -2546 -237 10154
rect 10449 10193 10543 10235
rect -150 10114 -90 10148
rect 10304 10114 10364 10148
rect -150 10088 10364 10114
rect -116 10065 10330 10088
rect -116 10015 48 10065
rect 10145 10015 10330 10065
rect -116 9970 10330 10015
rect -116 9936 27 9970
rect -116 -2341 -95 9936
rect -41 -2341 27 9936
rect 10175 9915 10330 9970
rect 10175 6151 10220 9915
rect 10272 6152 10330 9915
rect 10449 6344 10477 10193
rect 10534 6344 10543 10193
rect 12837 9463 12945 9473
rect 12837 9332 12850 9463
rect 12928 9332 12945 9463
rect 12837 9323 12945 9332
rect 12821 9011 12955 9026
rect 12821 8818 12834 9011
rect 12938 8818 12955 9011
rect 12821 8802 12955 8818
rect 11920 7236 12270 7248
rect 11920 7182 11945 7236
rect 12229 7182 12270 7236
rect 11920 7172 12270 7182
rect 10449 6313 10577 6344
rect 10449 6279 10615 6313
rect 11230 6279 11369 6313
rect 10449 6248 11369 6279
rect 10449 6186 11269 6248
rect 10272 6151 10364 6152
rect 10175 6067 10364 6151
rect 11086 6072 11156 6101
rect 11086 6067 11122 6072
rect 10175 6024 11122 6067
rect 10175 6008 11012 6024
rect 10175 5956 10226 6008
rect 10952 5956 11012 6008
rect 10175 5911 11012 5956
rect -116 -2346 27 -2341
rect 10966 -2346 11012 5911
rect -116 -2353 11012 -2346
rect 11068 -2353 11122 6024
rect -116 -2408 11122 -2353
rect -116 -2461 -4 -2408
rect 10961 -2461 11122 -2408
rect -116 -2466 11122 -2461
rect -116 -2475 11156 -2466
rect -150 -2501 11156 -2475
rect -150 -2535 -90 -2501
rect 11086 -2535 11156 -2501
rect -324 -2622 -237 -2546
rect 11241 -2594 11269 6186
rect 11326 -2594 11335 6248
rect 11241 -2622 11335 -2594
rect -324 -2651 11335 -2622
rect -324 -2686 -189 -2651
rect -358 -2691 -189 -2686
rect 11216 -2686 11335 -2651
rect 11216 -2691 11369 -2686
rect -358 -2712 11369 -2691
rect -358 -2746 -298 -2712
rect 11309 -2746 11369 -2712
<< viali >>
rect -216 10268 10415 10317
rect -312 -2546 -260 10154
rect 48 10015 10145 10065
rect -95 -2341 -41 9936
rect 10220 6151 10272 9915
rect 10477 6344 10534 10193
rect 12850 9332 12928 9463
rect 12834 8818 12938 9011
rect 11945 7182 12229 7236
rect 10226 5956 10952 6008
rect 11012 -2353 11068 6024
rect -4 -2461 10961 -2408
rect 11269 -2594 11326 6248
rect -189 -2691 11216 -2651
<< metal1 >>
rect -358 10317 10577 10357
rect -358 10268 -216 10317
rect 10415 10268 10577 10317
rect -358 10235 10577 10268
rect -358 10154 -237 10235
rect -358 -2546 -312 10154
rect -260 -2546 -237 10154
rect 10449 10193 10577 10235
rect -108 10065 10290 10085
rect -108 10015 48 10065
rect 10145 10015 10290 10065
rect -108 10002 10290 10015
rect -108 9936 -25 10002
rect 5161 9987 5347 10002
rect -108 -2341 -95 9936
rect -41 -2341 -25 9936
rect 10207 9915 10290 10002
rect 3896 6109 3942 6237
rect 10207 6151 10220 9915
rect 10272 6151 10290 9915
rect 10449 7635 10477 10193
rect 10377 7627 10477 7635
rect 10534 9689 10577 10193
rect 10534 9688 11709 9689
rect 10534 9554 11726 9688
rect 10534 7627 10577 9554
rect 10549 6801 10577 7627
rect 11626 7192 11726 9554
rect 11920 7236 12270 7248
rect 11610 6801 11758 7192
rect 11920 7182 11945 7236
rect 12229 7182 12270 7236
rect 12363 7196 12523 9684
rect 12861 9473 12913 9873
rect 12837 9463 12945 9473
rect 12837 9332 12850 9463
rect 12928 9332 12945 9463
rect 12837 9323 12945 9332
rect 12861 9026 12913 9323
rect 12821 9011 12955 9026
rect 12821 8818 12834 9011
rect 12938 8818 12955 9011
rect 12821 8802 12955 8818
rect 11920 7174 12028 7182
rect 12200 7174 12270 7182
rect 11920 7172 12270 7174
rect 12028 7168 12200 7172
rect 12322 7130 12572 7196
rect 12322 6873 12336 7130
rect 12558 6873 12572 7130
rect 12322 6854 12572 6873
rect 12600 7147 12657 7213
rect 13166 7199 13266 9686
rect 12600 7137 12742 7147
rect 12600 6861 12639 7137
rect 12731 6861 12742 7137
rect 12600 6851 12742 6861
rect 13136 6801 13284 7199
rect 10549 6794 13284 6801
rect 10549 6564 11031 6794
rect 11327 6564 13284 6794
rect 10549 6558 13284 6564
rect 10549 6344 10577 6558
rect 12047 6417 12053 6420
rect 10377 6331 10577 6344
rect 10746 6371 12053 6417
rect 10207 6142 10290 6151
rect 10746 6109 10792 6371
rect 12047 6368 12053 6371
rect 12225 6368 12231 6420
rect 11169 6248 11369 6261
rect 61 6063 10792 6109
rect 10866 6164 11104 6175
rect 61 4054 143 6063
rect 10866 6027 10875 6164
rect 10207 6008 10875 6027
rect 10207 5956 10226 6008
rect 10207 5944 10875 5956
rect 11093 5944 11104 6164
rect 10866 5935 11012 5944
rect 61 4008 664 4054
rect -108 -2390 -25 -2341
rect 10999 -2353 11012 5935
rect 11068 5935 11104 5944
rect 11068 -2353 11082 5935
rect 11341 5899 11369 6248
rect 11169 5891 11269 5899
rect 10999 -2390 11082 -2353
rect -108 -2408 11082 -2390
rect -108 -2461 -4 -2408
rect 10961 -2461 11082 -2408
rect -108 -2473 11082 -2461
rect -358 -2576 -237 -2546
rect -358 -2622 3257 -2576
rect 11241 -2594 11269 5891
rect 11326 -2594 11369 5899
rect 11448 5843 11680 5852
rect 11448 5746 11454 5843
rect 11673 5746 11680 5843
rect 11448 3913 11680 5746
rect 11448 3425 11455 3913
rect 11671 3425 11680 3913
rect 11448 3413 11680 3425
rect 11241 -2622 11369 -2594
rect -358 -2651 11369 -2622
rect -358 -2691 -189 -2651
rect 11216 -2691 11369 -2651
rect -358 -2746 11369 -2691
rect -355 -2799 3257 -2746
<< via1 >>
rect 10377 6344 10477 7627
rect 10477 6344 10534 7627
rect 10534 6344 10549 7627
rect 12028 7182 12200 7226
rect 12028 7174 12200 7182
rect 12336 6873 12558 7130
rect 12639 6861 12731 7137
rect 11031 6564 11327 6794
rect 12053 6368 12225 6420
rect 10875 6024 11093 6164
rect 10875 6008 11012 6024
rect 10875 5956 10952 6008
rect 10952 5956 11012 6008
rect 10875 5944 11012 5956
rect 11012 5944 11068 6024
rect 11068 5944 11093 6024
rect 11169 5899 11269 6248
rect 11269 5899 11326 6248
rect 11326 5899 11341 6248
rect 11454 5746 11673 5843
rect 11455 3425 11671 3913
<< metal2 >>
rect 5161 9987 5347 10085
rect 10353 7627 10576 7653
rect 10353 6344 10377 7627
rect 10549 6450 10576 7627
rect 12022 7223 12028 7226
rect 12014 7177 12028 7223
rect 12022 7174 12028 7177
rect 12200 7174 12206 7226
rect 11026 6794 11371 6802
rect 11026 6564 11031 6794
rect 11327 6564 11371 6794
rect 11026 6450 11371 6564
rect 10549 6344 11371 6450
rect 12096 6426 12161 7174
rect 12318 7130 12569 7143
rect 12318 6873 12336 7130
rect 12558 6873 12569 7130
rect 12053 6420 12225 6426
rect 12053 6362 12225 6368
rect 4961 6175 5147 6257
rect 10355 6248 11371 6344
rect 10355 6227 11169 6248
rect 9712 6164 11093 6175
rect 9712 6163 10875 6164
rect 9712 5949 9725 6163
rect 10824 5949 10875 6163
rect 9712 5944 10875 5949
rect 9712 5935 11093 5944
rect 4961 5914 5147 5935
rect 11129 5899 11169 6227
rect 11341 5899 11371 6248
rect 12318 6164 12569 6873
rect 12318 5948 12331 6164
rect 12552 5948 12569 6164
rect 12318 5936 12569 5948
rect 12630 7137 12741 7146
rect 12630 6861 12639 7137
rect 12731 6861 12741 7137
rect 11129 5865 11371 5899
rect 11113 4077 11371 5865
rect 12630 5849 12741 6861
rect 11437 5843 12741 5849
rect 11437 5746 11454 5843
rect 11673 5746 12741 5843
rect 11437 5738 12741 5746
rect 10640 3913 12121 3922
rect 10640 3425 11455 3913
rect 11671 3425 12121 3913
rect 10640 3417 12121 3425
rect -140 1871 198 1971
rect 10897 1738 11337 1838
rect -140 1636 198 1736
rect -140 1178 198 1278
<< via2 >>
rect 4961 5935 5147 6175
rect 9725 5949 10824 6163
rect 12331 5948 12552 6164
<< metal3 >>
rect 623 2142 723 7084
rect 1659 6114 1759 7545
rect 4954 6175 5158 6184
rect 835 6014 1759 6114
rect 2077 6160 4961 6175
rect 835 1343 935 6014
rect 2077 5948 2090 6160
rect 2488 5948 4961 6160
rect 2077 5935 4961 5948
rect 5147 6164 12571 6175
rect 5147 6163 12331 6164
rect 5147 5949 9725 6163
rect 10824 5949 12331 6163
rect 5147 5948 12331 5949
rect 12552 5948 12571 6164
rect 5147 5935 12571 5948
rect 4954 5927 5158 5935
<< via3 >>
rect 2090 5948 2488 6160
<< metal4 >>
rect 285 9775 1485 10036
rect 2570 9770 3770 10036
rect 285 6171 1485 6273
rect 2769 6216 6781 6936
rect 1685 6171 2501 6173
rect 285 6160 2501 6171
rect 285 5948 2090 6160
rect 2488 5948 2501 6160
rect 285 4660 2501 5948
rect 6061 5601 6781 6216
use cc_via2_3cut  cc_via2_3cut_0
timestamp 1717772055
transform 0 1 -639040 -1 0 518654
box 517199 639873 517310 640172
use cc_via2_3cut  cc_via2_3cut_1
timestamp 1717772055
transform 0 1 -639448 -1 0 519454
box 517199 639873 517310 640172
use comparator_bias  comparator_bias_0
timestamp 1747682096
transform -1 0 518254 0 1 -639855
box 508008 646042 518182 649916
use comparator_core_cload  comparator_core_cload_0
timestamp 1721179627
transform 1 0 -506133 0 1 -641069
box 506207 638825 517124 647001
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 1 11633 1 0 9302
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 13261 -1 0 9494
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 13261 -1 0 9686
box -66 -43 258 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 13261 -1 0 9302
box -66 -43 2178 1671
<< labels >>
flabel metal2 -140 1871 198 1971 0 FreeSans 1600 0 0 0 VINP
port 1 nsew
flabel metal2 -140 1636 198 1736 0 FreeSans 1600 0 0 0 VINM
port 0 nsew
flabel metal4 285 9775 1485 10036 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal4 2570 9770 3770 10036 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal2 11113 4077 11336 5865 0 FreeSans 1600 270 0 0 DVSS
port 6 nsew
flabel metal2 10902 3417 11337 3922 0 FreeSans 1600 0 0 0 DVDD
port 5 nsew
flabel metal2 10911 1738 11337 1838 0 FreeSans 1200 0 0 0 VOUT
port 7 nsew
flabel metal2 -140 1178 198 1278 0 FreeSans 1600 0 0 0 CLOAD
port 8 nsew
flabel metal1 12861 9704 12913 9873 0 FreeSans 320 90 0 0 ENA
port 9 nsew
<< end >>

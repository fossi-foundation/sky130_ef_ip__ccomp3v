magic
tech sky130A
magscale 1 2
timestamp 1747681386
<< error_s >>
rect 5080 -3224 5082 -3068
rect 5108 -3224 5110 -3096
<< dnwell >>
rect 2745 83 4814 1308
rect 2745 -267 4811 83
rect 289 -3321 4811 -267
<< nwell >>
rect 6286 1828 6496 2622
rect 2636 1464 3614 1522
rect 6286 1480 6428 1828
rect 2636 1462 4533 1464
rect 2636 1321 4671 1462
rect 2552 1270 4671 1321
rect 2552 132 2868 1270
rect 3740 1232 4671 1270
rect 3740 132 3958 1232
rect 2552 131 3958 132
rect 2552 -92 4670 131
rect 2552 -106 4946 -92
rect 138 -274 4946 -106
rect 138 -3276 306 -274
rect 4717 -3276 4946 -274
rect 138 -3444 4946 -3276
<< mvnsubdiff >>
rect 2772 1406 4737 1421
rect 2772 1367 2798 1406
rect 4568 1367 4737 1406
rect 2772 1349 4737 1367
rect 3822 1310 3880 1349
rect 3822 65 3831 1310
rect 3871 65 3880 1310
rect 3822 35 3880 65
rect 2852 15 4736 35
rect 2852 -24 2876 15
rect 4516 -24 4736 15
rect 2852 -36 4736 -24
rect 4818 -104 4880 -41
rect 4818 -3190 4828 -104
rect 4872 -3190 4880 -104
rect 4818 -3237 4880 -3190
<< mvnsubdiffcont >>
rect 2798 1367 4568 1406
rect 3831 65 3871 1310
rect 2876 -24 4516 15
rect 4828 -3190 4872 -104
<< locali >>
rect 3670 2989 4757 3004
rect 3670 2941 3729 2989
rect 4738 2941 4757 2989
rect 3670 2928 4757 2941
rect 3670 2880 3746 2928
rect 3670 1635 3684 2880
rect 3734 1635 3746 2880
rect 3670 1596 3746 1635
rect 4255 2880 4331 2928
rect 4255 1628 4272 2880
rect 4322 1628 4331 2880
rect 4255 1596 4331 1628
rect 4681 2880 4757 2928
rect 4681 1633 4690 2880
rect 4740 1633 4757 2880
rect 4681 1596 4757 1633
rect 4852 2982 6225 2998
rect 4852 2937 4872 2982
rect 6202 2937 6225 2982
rect 4852 2922 6225 2937
rect 4852 2880 4928 2922
rect 4852 1798 4865 2880
rect 4912 1798 4928 2880
rect 4852 1597 4928 1798
rect 6149 2878 6225 2922
rect 6149 1647 6166 2878
rect 6216 1647 6225 2878
rect 6556 2555 7051 2562
rect 6556 2505 6664 2555
rect 6811 2548 7051 2555
rect 6811 2505 6997 2548
rect 6556 2495 6997 2505
rect 6556 2481 6623 2495
rect 6556 2245 6566 2481
rect 6617 2245 6623 2481
rect 6556 1959 6623 2245
rect 6984 1963 6997 2495
rect 7041 1963 7051 2548
rect 6984 1959 7051 1963
rect 6556 1949 7051 1959
rect 6556 1902 6590 1949
rect 6951 1902 7051 1949
rect 6556 1893 7051 1902
rect 6556 1892 7042 1893
rect 6149 1597 6225 1647
rect 3670 1587 4758 1596
rect 3670 1535 3690 1587
rect 3975 1581 4604 1587
rect 3975 1535 4192 1581
rect 3670 1531 4192 1535
rect 4313 1536 4604 1581
rect 4745 1536 4758 1587
rect 4313 1531 4758 1536
rect 3670 1520 4758 1531
rect 4852 1581 6225 1597
rect 4852 1536 4992 1581
rect 6202 1536 6225 1581
rect 4852 1521 6225 1536
rect 4727 1421 6369 1425
rect 2770 1410 6369 1421
rect 2770 1406 2808 1410
rect 3244 1406 6369 1410
rect 2770 1367 2798 1406
rect 4568 1367 4748 1406
rect 2770 1359 4748 1367
rect 6345 1359 6369 1406
rect 2770 1349 6369 1359
rect 3824 1310 3880 1349
rect 2946 1180 3606 1197
rect 2946 1176 3449 1180
rect 2946 1137 2970 1176
rect 3270 1140 3449 1176
rect 3588 1140 3606 1180
rect 3270 1137 3606 1140
rect 2946 1121 3606 1137
rect 2946 1069 3022 1121
rect 2946 246 2965 1069
rect 3008 302 3022 1069
rect 3530 1066 3606 1121
rect 3530 302 3546 1066
rect 3008 285 3546 302
rect 3008 247 3056 285
rect 3507 247 3546 285
rect 3008 246 3546 247
rect 2946 243 3546 246
rect 3589 243 3606 1066
rect 2946 226 3606 243
rect 3824 65 3831 1310
rect 3871 1248 3880 1310
rect 3874 77 3880 1248
rect 4727 1312 4803 1349
rect 4036 1121 4541 1143
rect 4036 1118 4482 1121
rect 4036 295 4052 1118
rect 4095 1067 4482 1118
rect 4095 354 4112 1067
rect 4465 354 4482 1067
rect 4095 335 4482 354
rect 4095 298 4156 335
rect 4438 298 4482 335
rect 4525 298 4541 1121
rect 4095 295 4541 298
rect 4036 278 4541 295
rect 3871 65 3880 77
rect 3824 36 3880 65
rect 4727 54 4741 1312
rect 4788 54 4803 1312
rect 4727 36 4803 54
rect 2844 24 4803 36
rect 2844 15 2930 24
rect 4668 20 4803 24
rect 5510 1310 5586 1349
rect 5510 237 5529 1310
rect 5574 237 5586 1310
rect 5510 20 5586 237
rect 6293 1316 6369 1349
rect 6293 82 6309 1316
rect 6354 82 6369 1316
rect 6293 20 6369 82
rect 2844 -24 2876 15
rect 4668 14 6369 20
rect 4668 -17 4750 14
rect 4516 -24 4750 -17
rect 2844 -33 4750 -24
rect 6347 -33 6369 14
rect 2844 -36 6369 -33
rect 4727 -52 6369 -36
rect 4727 -56 6368 -52
rect 4818 -104 4880 -56
rect 384 -388 4626 -365
rect 384 -429 410 -388
rect 4605 -429 4626 -388
rect 384 -441 4626 -429
rect 384 -481 460 -441
rect 384 -1421 406 -481
rect 448 -1421 460 -481
rect 384 -1753 460 -1421
rect 3244 -479 3320 -441
rect 3244 -1525 3267 -479
rect 3308 -1525 3320 -479
rect 3244 -1753 3320 -1525
rect 4575 -491 4626 -441
rect 4575 -1753 4586 -491
rect 384 -1769 4586 -1753
rect 384 -1815 589 -1769
rect 4420 -1815 4586 -1769
rect 384 -1829 4586 -1815
rect 384 -2174 460 -1829
rect 384 -3096 405 -2174
rect 444 -3096 460 -2174
rect 384 -3136 460 -3096
rect 3244 -2036 3320 -1829
rect 3244 -3104 3264 -2036
rect 3301 -3104 3320 -2036
rect 3244 -3136 3320 -3104
rect 4575 -3099 4586 -1829
rect 4620 -3099 4626 -491
rect 4575 -3136 4626 -3099
rect 384 -3155 4626 -3136
rect 384 -3198 405 -3155
rect 4557 -3198 4626 -3155
rect 384 -3212 4626 -3198
rect 4818 -3190 4828 -104
rect 4875 -212 4880 -104
rect 4872 -355 4880 -212
rect 4875 -3164 4880 -355
rect 4872 -3190 4880 -3164
rect 4818 -3237 4880 -3190
rect 5019 -431 6299 -404
rect 5019 -471 5140 -431
rect 6275 -471 6299 -431
rect 5019 -480 6299 -471
rect 5019 -504 5095 -480
rect 5019 -1726 5041 -504
rect 5084 -1726 5095 -504
rect 5019 -1753 5095 -1726
rect 6223 -522 6299 -480
rect 6223 -1676 6242 -522
rect 6285 -1676 6299 -522
rect 6223 -1753 6299 -1676
rect 5019 -1829 6299 -1753
rect 5019 -1884 5095 -1829
rect 5019 -3075 5036 -1884
rect 5077 -3075 5095 -1884
rect 5019 -3136 5095 -3075
rect 6223 -1941 6299 -1829
rect 6223 -3082 6241 -1941
rect 6284 -3082 6299 -1941
rect 6223 -3136 6299 -3082
rect 5019 -3155 6299 -3136
rect 5019 -3198 5108 -3155
rect 6275 -3198 6299 -3155
rect 5019 -3212 6299 -3198
<< viali >>
rect 3729 2941 4738 2989
rect 3684 1635 3734 2880
rect 4272 1628 4322 2880
rect 4690 1633 4740 2880
rect 4872 2937 6202 2982
rect 4865 1798 4912 2880
rect 6166 1647 6216 2878
rect 6664 2505 6811 2555
rect 6566 2245 6617 2481
rect 6997 1963 7041 2548
rect 6590 1902 6951 1949
rect 3690 1535 3975 1587
rect 4192 1531 4313 1581
rect 4604 1536 4745 1587
rect 4992 1536 6202 1581
rect 2808 1406 3244 1410
rect 2808 1367 3244 1406
rect 4748 1359 6345 1406
rect 2970 1137 3270 1176
rect 3449 1140 3588 1180
rect 2965 246 3008 1069
rect 3056 247 3507 285
rect 3546 243 3589 1066
rect 3836 77 3871 1248
rect 3871 77 3874 1248
rect 4052 295 4095 1118
rect 4156 298 4438 335
rect 4482 298 4525 1121
rect 4741 54 4788 1312
rect 2930 15 4668 24
rect 5529 237 5574 1310
rect 6309 82 6354 1316
rect 2930 -17 4516 15
rect 4516 -17 4668 15
rect 4750 -33 6347 14
rect 410 -429 4605 -388
rect 406 -1421 448 -481
rect 3267 -1525 3308 -479
rect 589 -1815 4420 -1769
rect 405 -3096 444 -2174
rect 3264 -3104 3301 -2036
rect 4586 -3099 4620 -491
rect 405 -3198 4557 -3155
rect 4829 -212 4872 -104
rect 4872 -212 4875 -104
rect 4829 -3164 4872 -355
rect 4872 -3164 4875 -355
rect 5140 -471 6275 -431
rect 5041 -1726 5084 -504
rect 6242 -1676 6285 -522
rect 5036 -3075 5077 -1884
rect 6241 -3082 6284 -1941
rect 5108 -3198 6275 -3155
<< metal1 >>
rect 6804 3018 7004 3032
rect 3666 2989 4757 3004
rect 3666 2941 3729 2989
rect 4738 2941 4757 2989
rect 3666 2928 4757 2941
rect 3666 2880 3742 2928
rect 3666 1635 3684 2880
rect 3734 1635 3742 2880
rect 4258 2880 4334 2928
rect 3898 2818 3942 2824
rect 3776 2316 3862 2330
rect 3776 1768 3862 1780
rect 3898 1718 3928 2818
rect 4056 2816 4068 2822
rect 3958 2346 4042 2364
rect 3958 1800 4042 1816
rect 4070 1718 4102 2822
rect 4136 2472 4222 2486
rect 4136 1764 4222 1776
rect 3876 1672 4126 1718
rect 3666 1596 3742 1635
rect 3666 1587 3993 1596
rect 3666 1535 3690 1587
rect 3975 1535 3993 1587
rect 3666 1520 3993 1535
rect 2704 1410 3268 1424
rect 2704 1367 2808 1410
rect 3244 1367 3268 1410
rect 4070 1396 4110 1672
rect 4258 1628 4272 2880
rect 4322 1628 4334 2880
rect 4681 2880 4757 2928
rect 4258 1596 4334 1628
rect 4163 1581 4334 1596
rect 4163 1531 4192 1581
rect 4313 1531 4334 1581
rect 4163 1520 4334 1531
rect 2704 1349 3268 1367
rect 3334 1394 4209 1396
rect 4364 1394 4418 2748
rect 3334 1332 4418 1394
rect 4478 2120 4522 2826
rect 4562 2746 4646 2764
rect 4562 2200 4646 2216
rect 4478 2114 4530 2120
rect 4478 1748 4530 1754
rect 4478 1490 4522 1748
rect 4681 1633 4690 2880
rect 4740 1633 4757 2880
rect 4850 2982 6225 3000
rect 4850 2937 4872 2982
rect 6202 2937 6225 2982
rect 4850 2924 6225 2937
rect 4850 2880 4926 2924
rect 4850 1798 4865 2880
rect 4912 1798 4926 2880
rect 6149 2878 6225 2924
rect 4982 2746 5066 2764
rect 4982 2200 5066 2216
rect 4850 1764 4926 1798
rect 5130 1712 5174 2824
rect 5240 2472 5326 2482
rect 5240 1762 5326 1776
rect 5388 1712 5432 2824
rect 5498 2746 5582 2764
rect 5498 2200 5582 2216
rect 5646 1712 5690 2826
rect 5776 2482 5782 2484
rect 5816 2482 5822 2484
rect 5756 2472 5842 2482
rect 5756 1762 5842 1776
rect 5902 1712 5946 2822
rect 6014 2746 6098 2764
rect 6014 2198 6098 2216
rect 4681 1596 4757 1633
rect 4582 1587 4757 1596
rect 4582 1536 4604 1587
rect 4745 1536 4757 1587
rect 4786 1544 4800 1712
rect 4908 1664 6020 1712
rect 4908 1544 4920 1664
rect 6149 1647 6166 2878
rect 6216 1647 6225 2878
rect 6804 2654 6816 3018
rect 6990 2654 7004 3018
rect 6804 2640 7004 2654
rect 6556 2555 6834 2562
rect 6556 2548 6664 2555
rect 6556 2251 6563 2548
rect 6617 2505 6664 2548
rect 6811 2505 6834 2555
rect 6617 2496 6834 2505
rect 6556 2245 6566 2251
rect 6617 2245 6624 2496
rect 6556 2228 6624 2245
rect 6149 1597 6225 1647
rect 4962 1581 6225 1597
rect 4582 1520 4757 1536
rect 4962 1536 4992 1581
rect 6202 1536 6225 1581
rect 4962 1521 6225 1536
rect 6280 2124 6732 2192
rect 6280 1490 6324 2124
rect 6790 2075 6820 2404
rect 6882 2126 6926 2640
rect 6985 2548 7051 2562
rect 6985 2525 6997 2548
rect 7041 2525 7051 2548
rect 4478 1446 6324 1490
rect 6413 2045 6820 2075
rect 2946 1176 3286 1197
rect 2946 1137 2970 1176
rect 3270 1137 3286 1176
rect 2946 1121 3286 1137
rect 2946 1069 3022 1121
rect 2946 649 2965 1069
rect 3008 649 3022 1069
rect 3334 1040 3374 1332
rect 3824 1248 3881 1274
rect 3422 1180 3606 1197
rect 3422 1140 3449 1180
rect 3588 1140 3606 1180
rect 3422 1121 3606 1140
rect 3530 1066 3606 1121
rect 3154 994 3404 1040
rect 3088 954 3152 964
rect 3088 696 3152 706
rect 2946 289 2957 649
rect 3009 302 3022 649
rect 3182 392 3222 994
rect 3250 924 3306 940
rect 3250 458 3306 472
rect 3334 404 3374 994
rect 3408 956 3472 964
rect 3408 696 3472 708
rect 3530 651 3546 1066
rect 3589 651 3606 1066
rect 3530 302 3541 651
rect 3009 291 3541 302
rect 3594 291 3606 651
rect 3009 289 3546 291
rect 2946 246 2965 289
rect 3008 285 3546 289
rect 3008 247 3056 285
rect 3507 247 3546 285
rect 3008 246 3546 247
rect 2946 243 3546 246
rect 3589 243 3606 291
rect 2946 226 3606 243
rect 3824 77 3836 1248
rect 3874 77 3881 1248
rect 4035 1118 4111 1142
rect 4035 686 4052 1118
rect 4095 686 4111 1118
rect 4035 300 4046 686
rect 4099 354 4111 686
rect 4149 514 4209 1332
rect 4478 1254 4522 1446
rect 4273 1218 4522 1254
rect 4725 1410 6372 1413
rect 4725 1406 4749 1410
rect 6342 1406 6372 1410
rect 4725 1359 4748 1406
rect 6345 1359 6372 1406
rect 4725 1346 4749 1359
rect 6342 1346 6372 1359
rect 4725 1337 6372 1346
rect 4725 1312 4801 1337
rect 4725 1302 4741 1312
rect 4788 1302 4801 1312
rect 4273 452 4309 1218
rect 4465 1121 4541 1143
rect 4361 898 4417 908
rect 4361 512 4417 526
rect 4465 354 4482 1121
rect 4099 335 4482 354
rect 4099 300 4156 335
rect 4035 295 4052 300
rect 4095 298 4156 300
rect 4438 298 4482 335
rect 4525 298 4541 1121
rect 4095 295 4541 298
rect 4035 278 4541 295
rect 4725 794 4740 1302
rect 4795 794 4801 1302
rect 5511 1310 5587 1337
rect 5511 1295 5529 1310
rect 5574 1295 5587 1310
rect 3824 36 3881 77
rect 4725 54 4741 794
rect 4788 54 4801 794
rect 4864 1168 4940 1186
rect 4864 788 4940 802
rect 5004 144 5048 1258
rect 5112 624 5198 640
rect 5112 196 5198 210
rect 5258 144 5302 1244
rect 5380 1168 5456 1186
rect 5380 788 5456 802
rect 5511 787 5523 1295
rect 5578 787 5587 1295
rect 6293 1316 6369 1337
rect 6293 1304 6309 1316
rect 6354 1304 6369 1316
rect 5648 1168 5724 1186
rect 5648 788 5724 802
rect 5511 237 5529 787
rect 5574 237 5587 787
rect 5511 213 5587 237
rect 4928 142 5386 144
rect 5790 142 5834 1248
rect 5896 620 5982 636
rect 5896 142 5982 206
rect 6042 142 6086 1248
rect 6164 1168 6240 1186
rect 6164 788 6240 802
rect 6293 796 6303 1304
rect 6358 796 6369 1304
rect 4928 96 6170 142
rect 5380 94 6170 96
rect 4725 36 4801 54
rect 2706 24 4801 36
rect 6293 82 6309 796
rect 6354 82 6369 796
rect 6293 24 6369 82
rect 2706 -17 2930 24
rect 4668 14 6369 24
rect 4668 -17 4750 14
rect 2706 -33 4750 -17
rect 6347 -33 6369 14
rect 2706 -37 6369 -33
rect 4725 -52 6369 -37
rect 4806 -104 4892 -52
rect 4806 -212 4829 -104
rect 4875 -212 4892 -104
rect 4806 -234 4892 -212
rect 4806 -355 4892 -334
rect 386 -368 4618 -364
rect 386 -377 4626 -368
rect 386 -430 392 -377
rect 4520 -388 4626 -377
rect 4605 -429 4626 -388
rect 4520 -430 4626 -429
rect 386 -440 4626 -430
rect 386 -481 462 -440
rect 386 -526 406 -481
rect 448 -526 462 -481
rect 386 -1420 399 -526
rect 454 -1420 462 -526
rect 3244 -479 3320 -440
rect 528 -642 596 -610
rect 528 -1044 596 -1016
rect 386 -1421 406 -1420
rect 448 -1421 462 -1420
rect 386 -1442 462 -1421
rect 228 -1515 490 -1506
rect 228 -1699 229 -1515
rect 290 -1630 490 -1515
rect 668 -1630 708 -536
rect 792 -1166 852 -1114
rect 792 -1578 852 -1560
rect 926 -1630 966 -536
rect 1044 -642 1112 -610
rect 1044 -1044 1112 -1016
rect 1184 -1630 1224 -536
rect 1308 -1166 1368 -1114
rect 1308 -1578 1368 -1560
rect 1442 -1630 1482 -536
rect 1560 -642 1628 -610
rect 1560 -1044 1628 -1016
rect 1700 -1630 1740 -536
rect 1824 -1166 1884 -1114
rect 1824 -1578 1884 -1560
rect 1958 -1630 1998 -536
rect 2076 -642 2144 -610
rect 2076 -1044 2144 -1016
rect 2216 -1630 2256 -536
rect 2340 -1166 2400 -1114
rect 2340 -1578 2400 -1560
rect 2474 -1630 2514 -536
rect 2592 -642 2660 -610
rect 2592 -1044 2660 -1016
rect 2732 -1630 2772 -536
rect 2856 -1166 2916 -1114
rect 2856 -1578 2916 -1560
rect 2990 -1630 3030 -536
rect 3108 -642 3176 -610
rect 3108 -1044 3176 -1016
rect 3244 -1525 3267 -479
rect 3308 -1525 3320 -479
rect 4575 -491 4626 -440
rect 3244 -1546 3320 -1525
rect 3398 -1166 3458 -1114
rect 3398 -1578 3458 -1560
rect 3532 -1630 3572 -540
rect 3648 -642 3720 -612
rect 3648 -1034 3720 -1016
rect 3798 -1630 3838 -534
rect 3914 -1166 3974 -1114
rect 3914 -1578 3974 -1560
rect 4054 -1630 4094 -536
rect 4164 -642 4236 -612
rect 4164 -1034 4236 -1016
rect 4310 -1630 4350 -536
rect 4575 -643 4586 -491
rect 4430 -1166 4490 -1114
rect 4430 -1578 4490 -1560
rect 290 -1682 4350 -1630
rect 290 -1699 490 -1682
rect 228 -1706 490 -1699
rect 228 -1707 290 -1706
rect 556 -1764 4444 -1753
rect 556 -1769 618 -1764
rect 4413 -1769 4444 -1764
rect 556 -1815 589 -1769
rect 4420 -1815 4444 -1769
rect 556 -1819 618 -1815
rect 4413 -1819 4444 -1815
rect 556 -1829 4444 -1819
rect 229 -1866 291 -1865
rect 229 -1873 490 -1866
rect 229 -2057 230 -1873
rect 291 -1878 490 -1873
rect 291 -1930 4344 -1878
rect 291 -2057 490 -1930
rect 229 -2066 490 -2057
rect 528 -1994 596 -1984
rect 384 -2174 460 -2142
rect 384 -2187 405 -2174
rect 444 -2187 460 -2174
rect 384 -2725 392 -2187
rect 446 -2725 460 -2187
rect 528 -2416 596 -2368
rect 384 -3096 405 -2725
rect 444 -3096 460 -2725
rect 666 -3046 706 -1930
rect 790 -2520 850 -2488
rect 790 -2970 850 -2910
rect 924 -3046 964 -1930
rect 1044 -1994 1112 -1984
rect 1044 -2416 1112 -2368
rect 1182 -3046 1222 -1930
rect 1306 -2520 1366 -2490
rect 1306 -2970 1366 -2910
rect 1440 -3046 1480 -1930
rect 1560 -1994 1628 -1984
rect 1560 -2416 1628 -2368
rect 1698 -3046 1738 -1930
rect 1822 -2520 1882 -2496
rect 1822 -2970 1882 -2910
rect 1956 -3046 1996 -1930
rect 2076 -1994 2144 -1984
rect 2076 -2416 2144 -2368
rect 2214 -3046 2254 -1930
rect 2338 -2520 2398 -2500
rect 2338 -2970 2398 -2910
rect 2472 -3046 2512 -1930
rect 2592 -1994 2660 -1984
rect 2592 -2416 2660 -2368
rect 2730 -3046 2770 -1930
rect 2854 -2520 2914 -2492
rect 2854 -2970 2914 -2910
rect 2988 -3046 3028 -1930
rect 3108 -1994 3176 -1984
rect 3108 -2416 3176 -2368
rect 3251 -2036 3327 -2015
rect 384 -3136 460 -3096
rect 3251 -3104 3264 -2036
rect 3301 -3104 3327 -2036
rect 3396 -2520 3456 -2478
rect 3396 -2970 3456 -2910
rect 3532 -3048 3572 -1930
rect 3650 -1994 3722 -1982
rect 3650 -2404 3722 -2368
rect 3792 -3046 3832 -1930
rect 3912 -2520 3972 -2478
rect 3912 -2970 3972 -2910
rect 4048 -3050 4088 -1930
rect 4166 -1994 4238 -1982
rect 4166 -2404 4238 -2368
rect 4304 -3044 4344 -1930
rect 4572 -2368 4586 -643
rect 4620 -643 4626 -491
rect 4620 -665 4660 -643
rect 4647 -2344 4660 -665
rect 4428 -2520 4488 -2478
rect 4428 -2970 4488 -2910
rect 3251 -3136 3327 -3104
rect 4575 -3099 4586 -2368
rect 4620 -2368 4660 -2344
rect 4620 -3099 4626 -2368
rect 4575 -3136 4626 -3099
rect 384 -3143 4626 -3136
rect 384 -3155 424 -3143
rect 384 -3198 405 -3155
rect 4557 -3198 4626 -3143
rect 384 -3212 4626 -3198
rect 4806 -3164 4829 -355
rect 4875 -3164 4892 -355
rect 4806 -3260 4892 -3164
rect 5027 -424 6300 -408
rect 5027 -476 5056 -424
rect 6272 -431 6300 -424
rect 6275 -471 6300 -431
rect 6272 -476 6300 -471
rect 5027 -484 6300 -476
rect 5027 -504 5103 -484
rect 5027 -1837 5041 -504
rect 5084 -513 5103 -504
rect 5095 -1837 5103 -513
rect 6224 -522 6300 -484
rect 5166 -642 5234 -634
rect 5166 -1024 5234 -1016
rect 5027 -1884 5103 -1837
rect 5027 -3075 5036 -1884
rect 5077 -3075 5103 -1884
rect 5398 -1760 5484 -570
rect 5606 -1158 5722 -1148
rect 5606 -1576 5614 -1158
rect 5702 -1576 5722 -1158
rect 5606 -1586 5722 -1576
rect 5850 -1760 5936 -574
rect 6082 -642 6150 -634
rect 6082 -1024 6150 -1016
rect 6224 -1683 6238 -522
rect 6292 -1683 6300 -522
rect 6413 -1054 6443 2045
rect 6985 1958 6991 2525
rect 6556 1949 6991 1958
rect 6556 1902 6590 1949
rect 6951 1926 6991 1949
rect 6951 1902 7051 1926
rect 6556 1894 7051 1902
rect 6965 1892 7051 1894
rect 6413 -1254 6506 -1054
rect 6445 -1386 6475 -1254
rect 6445 -1398 6522 -1386
rect 6445 -1628 6468 -1398
rect 6445 -1640 6522 -1628
rect 6445 -1641 6475 -1640
rect 6224 -1697 6300 -1683
rect 6504 -1760 6704 -1698
rect 5398 -1828 6704 -1760
rect 5170 -1994 5234 -1980
rect 5170 -2388 5234 -2368
rect 5398 -3038 5484 -1828
rect 5608 -2548 5714 -2536
rect 5608 -2956 5620 -2548
rect 5704 -2956 5714 -2548
rect 5608 -2971 5714 -2956
rect 5850 -3042 5936 -1828
rect 6504 -1898 6704 -1828
rect 6223 -1921 6299 -1909
rect 6086 -1994 6150 -1980
rect 6086 -2388 6150 -2368
rect 6223 -2723 6238 -1921
rect 6293 -2723 6299 -1921
rect 5027 -3136 5103 -3075
rect 6223 -3082 6241 -2723
rect 6284 -3082 6299 -2723
rect 6223 -3136 6299 -3082
rect 5027 -3143 6299 -3136
rect 5027 -3198 5108 -3143
rect 6275 -3198 6299 -3143
rect 5027 -3212 6299 -3198
<< via1 >>
rect 3776 1780 3862 2316
rect 3958 1816 4042 2346
rect 4136 1776 4222 2472
rect 4562 2216 4646 2746
rect 4478 1754 4530 2114
rect 4982 2216 5066 2746
rect 5240 1776 5326 2472
rect 5498 2216 5582 2746
rect 5756 1776 5842 2472
rect 6014 2216 6098 2746
rect 4800 1544 4908 1712
rect 6816 2654 6990 3018
rect 6563 2481 6617 2548
rect 6563 2251 6566 2481
rect 6566 2251 6617 2481
rect 3088 706 3152 954
rect 2957 289 2965 649
rect 2965 289 3008 649
rect 3008 289 3009 649
rect 3250 472 3306 924
rect 3408 708 3472 956
rect 3541 291 3546 651
rect 3546 291 3589 651
rect 3589 291 3594 651
rect 4046 300 4052 686
rect 4052 300 4095 686
rect 4095 300 4099 686
rect 4749 1406 6342 1410
rect 4749 1359 6342 1406
rect 4749 1346 6342 1359
rect 4361 526 4417 898
rect 4740 794 4741 1302
rect 4741 794 4788 1302
rect 4788 794 4795 1302
rect 4864 802 4940 1168
rect 5112 210 5198 624
rect 5380 802 5456 1168
rect 5523 787 5529 1295
rect 5529 787 5574 1295
rect 5574 787 5578 1295
rect 5648 802 5724 1168
rect 5896 206 5982 620
rect 6164 802 6240 1168
rect 6303 796 6309 1304
rect 6309 796 6354 1304
rect 6354 796 6358 1304
rect 392 -388 4520 -377
rect 392 -429 410 -388
rect 410 -429 4520 -388
rect 392 -430 4520 -429
rect 399 -1420 406 -526
rect 406 -1420 448 -526
rect 448 -1420 454 -526
rect 528 -1016 596 -642
rect 229 -1699 290 -1515
rect 792 -1560 852 -1166
rect 1044 -1016 1112 -642
rect 1308 -1560 1368 -1166
rect 1560 -1016 1628 -642
rect 1824 -1560 1884 -1166
rect 2076 -1016 2144 -642
rect 2340 -1560 2400 -1166
rect 2592 -1016 2660 -642
rect 2856 -1560 2916 -1166
rect 3108 -1016 3176 -642
rect 3398 -1560 3458 -1166
rect 3648 -1016 3720 -642
rect 3914 -1560 3974 -1166
rect 4164 -1016 4236 -642
rect 4430 -1560 4490 -1166
rect 618 -1769 4413 -1764
rect 618 -1815 4413 -1769
rect 618 -1819 4413 -1815
rect 230 -2057 291 -1873
rect 392 -2725 405 -2187
rect 405 -2725 444 -2187
rect 444 -2725 446 -2187
rect 528 -2368 596 -1994
rect 790 -2910 850 -2520
rect 1044 -2368 1112 -1994
rect 1306 -2910 1366 -2520
rect 1560 -2368 1628 -1994
rect 1822 -2910 1882 -2520
rect 2076 -2368 2144 -1994
rect 2338 -2910 2398 -2520
rect 2592 -2368 2660 -1994
rect 2854 -2910 2914 -2520
rect 3108 -2368 3176 -1994
rect 3396 -2910 3456 -2520
rect 3650 -2368 3722 -1994
rect 3912 -2910 3972 -2520
rect 4166 -2368 4238 -1994
rect 4592 -2344 4620 -665
rect 4620 -2344 4647 -665
rect 4428 -2910 4488 -2520
rect 424 -3155 4557 -3143
rect 424 -3196 4557 -3155
rect 5056 -431 6272 -424
rect 5056 -471 5140 -431
rect 5140 -471 6272 -431
rect 5056 -476 6272 -471
rect 5041 -1726 5084 -513
rect 5084 -1726 5095 -513
rect 5041 -1837 5095 -1726
rect 5166 -1016 5234 -642
rect 5614 -1576 5702 -1158
rect 6082 -1016 6150 -642
rect 6238 -1676 6242 -522
rect 6242 -1676 6285 -522
rect 6285 -1676 6292 -522
rect 6238 -1683 6292 -1676
rect 6991 1963 6997 2525
rect 6997 1963 7041 2525
rect 7041 1963 7051 2525
rect 6991 1926 7051 1963
rect 6468 -1628 6522 -1398
rect 5170 -2368 5234 -1994
rect 5620 -2956 5704 -2548
rect 6086 -2368 6150 -1994
rect 6238 -1941 6293 -1921
rect 6238 -2723 6241 -1941
rect 6241 -2723 6284 -1941
rect 6284 -2723 6293 -1941
rect 5108 -3155 6275 -3143
rect 5108 -3196 6275 -3155
<< metal2 >>
rect 2664 3018 7124 3348
rect 2664 2746 6816 3018
rect 2664 2640 4562 2746
rect 2664 2368 4042 2574
rect 3958 2346 4042 2368
rect 3772 2316 3866 2334
rect 3772 1780 3776 2316
rect 3862 1780 3866 2316
rect 3958 1800 4042 1816
rect 4130 2472 4224 2490
rect 3772 1486 3866 1780
rect 3742 1484 3866 1486
rect 4130 1776 4136 2472
rect 4222 1776 4224 2472
rect 4646 2640 4982 2746
rect 4562 2200 4646 2216
rect 5066 2640 5498 2746
rect 4982 2200 5066 2216
rect 5240 2472 5326 2482
rect 4130 1484 4224 1776
rect 4452 1754 4478 2114
rect 4530 1776 5240 2114
rect 5582 2640 6014 2746
rect 5498 2200 5582 2216
rect 5756 2472 5842 2482
rect 5326 2110 5756 2114
rect 5326 1776 5328 2110
rect 4530 1762 5328 1776
rect 5456 1776 5756 2110
rect 6098 2654 6816 2746
rect 6990 2654 7124 3018
rect 6098 2640 7124 2654
rect 6014 2198 6098 2216
rect 6252 2548 6631 2640
rect 6252 2251 6563 2548
rect 6617 2251 6631 2548
rect 5842 1776 6098 2114
rect 5456 1762 6098 1776
rect 4530 1754 6098 1762
rect 6252 1895 6631 2251
rect 6974 2525 7078 2640
rect 6974 1926 6991 2525
rect 7051 1926 7078 2525
rect 4786 1618 4800 1712
rect 3022 1198 4224 1484
rect 4596 1544 4800 1618
rect 4908 1544 4920 1712
rect 3070 954 3174 1198
rect 3070 706 3088 954
rect 3152 706 3174 954
rect 3386 956 3490 1198
rect 3070 694 3174 706
rect 3250 924 3306 940
rect 2676 649 3250 658
rect 2676 289 2957 649
rect 3009 472 3250 649
rect 3386 708 3408 956
rect 3472 708 3490 956
rect 4361 898 4417 908
rect 3386 696 3490 708
rect 4029 686 4361 708
rect 3306 651 3596 658
rect 3306 472 3541 651
rect 3009 291 3541 472
rect 3594 291 3596 651
rect 3009 289 3596 291
rect 2676 276 3596 289
rect 4029 300 4046 686
rect 4099 526 4361 686
rect 4417 526 4445 708
rect 4099 300 4445 526
rect 4029 195 4445 300
rect 4029 68 4041 195
rect 4437 68 4445 195
rect 4029 58 4445 68
rect 4596 28 4670 1544
rect 6252 1460 6466 1895
rect 6974 1868 7078 1926
rect 4730 1410 6466 1460
rect 4730 1346 4749 1410
rect 6342 1346 6466 1410
rect 4730 1304 6466 1346
rect 4730 1302 6303 1304
rect 4730 794 4740 1302
rect 4795 1295 6303 1302
rect 4795 1168 5523 1295
rect 4795 802 4864 1168
rect 4940 802 5380 1168
rect 5456 802 5523 1168
rect 4795 794 5523 802
rect 4730 787 5523 794
rect 5578 1168 6303 1295
rect 5578 802 5648 1168
rect 5724 802 6164 1168
rect 6240 802 6303 1168
rect 5578 796 6303 802
rect 6358 796 6466 1304
rect 5578 787 6466 796
rect 4730 782 6466 787
rect 5105 624 5223 649
rect 5105 210 5112 624
rect 5198 210 5223 624
rect 5105 28 5223 210
rect 2667 26 5223 28
rect 2667 -86 2696 26
rect 3064 -86 5223 26
rect 2667 -90 5223 -86
rect 5875 620 5993 641
rect 5875 206 5896 620
rect 5982 206 5993 620
rect 5875 -166 5993 206
rect 2922 -168 5993 -166
rect 2922 -280 2952 -168
rect 3320 -280 5993 -168
rect 2922 -284 5993 -280
rect 4996 -354 5115 -353
rect 334 -377 4618 -354
rect 334 -430 392 -377
rect 4520 -430 4618 -377
rect 334 -482 4618 -430
rect 4996 -367 6406 -354
rect 334 -526 462 -482
rect 334 -1420 399 -526
rect 454 -1420 462 -526
rect 509 -1016 528 -642
rect 596 -1016 1044 -642
rect 1112 -1016 1560 -642
rect 1628 -1016 2076 -642
rect 2144 -1016 2592 -642
rect 2660 -1016 2696 -642
rect 2810 -1016 3108 -642
rect 3176 -1016 3212 -642
rect 3354 -1016 3648 -642
rect 3720 -1016 4164 -642
rect 4236 -665 4930 -642
rect 4236 -1016 4592 -665
rect 69 -1515 290 -1506
rect 69 -1699 229 -1515
rect 69 -1707 290 -1699
rect 334 -1718 462 -1420
rect 588 -1560 792 -1166
rect 852 -1560 1308 -1166
rect 1368 -1560 1824 -1166
rect 1884 -1560 2340 -1166
rect 2400 -1560 2856 -1166
rect 2916 -1560 3398 -1166
rect 3458 -1560 3914 -1166
rect 3974 -1560 4430 -1166
rect 4490 -1560 4502 -1166
rect 334 -1764 4438 -1718
rect 334 -1819 618 -1764
rect 4413 -1819 4438 -1764
rect 334 -1844 4438 -1819
rect 70 -1873 291 -1865
rect 70 -2057 230 -1873
rect 70 -2066 291 -2057
rect 334 -2187 462 -1844
rect 4532 -1994 4592 -1016
rect 334 -2725 392 -2187
rect 446 -2725 462 -2187
rect 515 -2368 528 -1994
rect 596 -2368 1044 -1994
rect 1112 -2368 1560 -1994
rect 1628 -2368 2076 -1994
rect 2144 -2368 2592 -1994
rect 2660 -2366 2954 -1994
rect 3068 -2366 3108 -1994
rect 2660 -2368 3108 -2366
rect 3176 -2368 3214 -1994
rect 3356 -2368 3650 -1994
rect 3722 -2368 4166 -1994
rect 4238 -2344 4592 -1994
rect 4647 -1994 4930 -665
rect 4996 -1000 5008 -367
rect 5103 -424 6406 -367
rect 6272 -476 6406 -424
rect 5103 -482 6406 -476
rect 5103 -1000 5115 -482
rect 6213 -522 6406 -482
rect 4996 -1837 5041 -1000
rect 5095 -1837 5115 -1000
rect 5158 -1016 5166 -642
rect 5234 -646 6082 -642
rect 5234 -1008 5330 -646
rect 5456 -1008 6082 -646
rect 5234 -1016 6082 -1008
rect 6150 -1016 6162 -642
rect 6213 -1148 6238 -522
rect 4996 -1910 5115 -1837
rect 5200 -1158 6238 -1148
rect 5200 -1576 5614 -1158
rect 5702 -1576 6238 -1158
rect 5200 -1683 6238 -1576
rect 6292 -1683 6406 -522
rect 5200 -1844 6406 -1683
rect 6468 -1398 6522 -1386
rect 6468 -1750 6522 -1628
rect 6206 -1921 6406 -1844
rect 4647 -2344 5170 -1994
rect 4238 -2368 5170 -2344
rect 5234 -2368 6086 -1994
rect 6150 -2368 6156 -1994
rect 334 -3096 462 -2725
rect 548 -2910 790 -2520
rect 850 -2910 1306 -2520
rect 1366 -2910 1822 -2520
rect 1882 -2910 2338 -2520
rect 2398 -2910 2854 -2520
rect 2914 -2910 3396 -2520
rect 3456 -2910 3912 -2520
rect 3972 -2910 4428 -2520
rect 4488 -2910 4526 -2520
rect 548 -2914 4526 -2910
rect 334 -3143 4557 -3096
rect 334 -3196 424 -3143
rect 334 -3224 4557 -3196
rect 4679 -3224 5082 -2516
rect 6206 -2536 6238 -1921
rect 5146 -2548 6238 -2536
rect 5146 -2956 5620 -2548
rect 5704 -2723 6238 -2548
rect 6293 -2723 6406 -1921
rect 5704 -2956 6406 -2723
rect 5146 -3096 6406 -2956
rect 5108 -3143 6406 -3096
rect 6275 -3196 6406 -3143
rect 5108 -3224 6406 -3196
<< via2 >>
rect 5328 1762 5456 2110
rect 4041 68 4437 195
rect 2696 -86 3064 26
rect 2952 -280 3320 -168
rect 2696 -1016 2810 -642
rect 2954 -2366 3068 -1994
rect 5008 -424 5103 -367
rect 5008 -476 5056 -424
rect 5056 -476 5103 -424
rect 5008 -513 5103 -476
rect 5008 -1000 5041 -513
rect 5041 -1000 5095 -513
rect 5095 -1000 5103 -513
rect 5330 -1008 5456 -646
<< metal3 >>
rect 5322 2110 5462 2120
rect 5322 1762 5328 2110
rect 5456 1762 5462 2110
rect 4029 195 4446 205
rect 4029 68 4041 195
rect 4437 68 4446 195
rect 2688 26 3074 32
rect 2688 -86 2696 26
rect 3064 -86 3074 26
rect 2688 -94 3074 -86
rect 4029 -60 4446 68
rect 2688 -642 2818 -94
rect 2942 -168 3328 -162
rect 2942 -280 2952 -168
rect 3320 -280 3328 -168
rect 4029 -185 5115 -60
rect 2942 -288 3328 -280
rect 2688 -1016 2696 -642
rect 2810 -1016 2818 -642
rect 2688 -2930 2818 -1016
rect 2946 -1994 3076 -288
rect 4990 -367 5115 -185
rect 4990 -1000 5008 -367
rect 5103 -1000 5115 -367
rect 4990 -1013 5115 -1000
rect 5322 -646 5462 1762
rect 5322 -1008 5330 -646
rect 5456 -1008 5462 -646
rect 5322 -1027 5462 -1008
rect 2946 -2366 2954 -1994
rect 3068 -2366 3076 -1994
rect 2946 -2927 3076 -2366
use sky130_fd_pr__nfet_05v0_nvt_N7RQJ6  sky130_fd_pr__nfet_05v0_nvt_N7RQJ6_0 paramcells
timestamp 1731019923
transform -1 0 1853 0 1 -1082
box -1497 -758 1497 758
use sky130_fd_pr__nfet_g5v0d10v5_R6PXNO  sky130_fd_pr__nfet_g5v0d10v5_R6PXNO_0 paramcells
timestamp 1731019923
transform -1 0 3943 0 1 -1082
box -723 -758 723 758
use sky130_fd_pr__pfet_g5v0d10v5_5FCQ7L  sky130_fd_pr__pfet_g5v0d10v5_5FCQ7L_0 paramcells
timestamp 1731019923
transform -1 0 4001 0 -1 2259
box -387 -797 387 797
use sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ  sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ_0 paramcells
timestamp 1731019923
transform 1 0 5157 0 1 683
box -487 -797 487 797
use sky130_fd_pr__nfet_g5v0d10v5_R6PXNO  XM2
timestamp 1731019923
transform -1 0 3943 0 1 -2468
box -723 -758 723 758
use sky130_fd_pr__nfet_g5v0d10v5_25MXQV  XM3 paramcells
timestamp 1731019923
transform -1 0 5661 0 1 -2468
box -665 -758 665 758
use sky130_fd_pr__nfet_05v0_nvt_N7RQJ6  XM5
timestamp 1731019923
transform -1 0 1853 0 1 -2468
box -1497 -758 1497 758
use sky130_fd_pr__pfet_g5v0d10v5_3P3PJP  XM8 paramcells
timestamp 1731019923
transform 1 0 6804 0 1 2225
box -308 -397 308 397
use sky130_fd_pr__pfet_g5v0d10v5_CBUN3Q  XM9 paramcells
timestamp 1731019923
transform -1 0 5541 0 1 2259
box -745 -797 745 797
use sky130_fd_pr__nfet_g5v0d10v5_D5V3WB  XM10 paramcells
timestamp 1731019923
transform -1 0 5661 0 1 -1102
box -665 -738 665 738
use sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ  XM12
timestamp 1731019923
transform 1 0 5941 0 1 683
box -487 -797 487 797
use sky130_fd_pr__pfet_g5v0d10v5_6THU7R  XM19 paramcells
timestamp 1731019923
transform -1 0 4506 0 -1 2259
box -308 -797 308 797
use sky130_fd_pr__nfet_g5v0d10v5_VR3TSB  XM20 paramcells
timestamp 1731019923
transform -1 0 4289 0 -1 712
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_TEGW2X  XM22 paramcells
timestamp 1731019923
transform -1 0 3279 0 -1 712
box -357 -508 357 508
<< labels >>
flabel metal2 2674 2372 2874 2572 0 FreeSans 256 0 0 0 DVDD
port 6 nsew
flabel metal2 2676 366 2876 566 0 FreeSans 256 0 0 0 DVSS
port 8 nsew
flabel metal2 3026 2852 3226 3052 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal2 6108 -2956 6308 -2756 0 FreeSans 256 180 0 0 VSS
port 2 nsew
flabel metal1 6504 -1898 6704 -1698 0 FreeSans 256 0 0 0 VBN
port 1 nsew
flabel metal1 6413 -1254 6506 -1054 0 FreeSans 256 0 0 0 ena3v3
port 7 nsew
flabel metal1 290 -2066 490 -1866 0 FreeSans 256 0 0 0 VINM
port 5 nsew
flabel metal1 290 -1706 490 -1506 0 FreeSans 256 0 0 0 VINP
port 3 nsew
flabel metal2 3046 1252 3246 1452 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
<< end >>

** sch_path: /home/tim/gits/sky130_ef_ip__ccomp3v/xschem/sky130_ef_ip__scomp3v.sch
.subckt sky130_ef_ip__scomp3v VOUT DVDD DVSS VDD VSS VINP VINM ENA
*.PININFO VDD:I VOUT:O VSS:I VINP:I VINM:I DVDD:I DVSS:I ENA:I
x3 ENA DVDD DVSS DVSS VDD VDD ena3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x1 VDD VBN VSS VINP VOUT VINM DVDD ena3v3 DVSS comparator_high_gain
x2 VDD VSS VBN ena3v3 scomp_bias
x4 ENA DVSS DVSS VDD VDD sky130_fd_sc_hvl__diode_2
.ends

* expanding   symbol:  comparator_high_gain.sym # of pins=9
** sym_path: /home/tim/gits/sky130_ef_ip__ccomp3v/xschem/comparator_high_gain.sym
** sch_path: /home/tim/gits/sky130_ef_ip__ccomp3v/xschem/comparator_high_gain.sch
.subckt comparator_high_gain VDD VBN VSS VINP VOUT VINM DVDD ena3v3 DVSS
*.PININFO VINP:I VINM:I VBN:I VDD:B VSS:B VOUT:O DVDD:B ena3v3:I DVSS:B
XM3 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM19 net2 VOUTANALOG VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM20 net2 VOUTANALOG VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM21 VOUT net2 DVDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM22 VOUT net2 DVSS DVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM1 net4 VINM net1 net1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM4 net6 VINM net4 net1 sky130_fd_pr__nfet_05v0_nvt L=1 W=5 nf=1 m=10
XM5 net5 VINP net3 net1 sky130_fd_pr__nfet_05v0_nvt L=1 W=5 nf=1 m=10
XM8 VOUTANALOG ena3v3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTANALOG net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=2 m=2
XM10 VOUTANALOG VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4.8 nf=1 m=2
XM11 net8 net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
XM12 net7 net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
Vmeas net8 net6 0
.save i(vmeas)
Vmeas1 net7 net5 0
.save i(vmeas1)
.ends


* expanding   symbol:  scomp_bias.sym # of pins=4
** sym_path: /home/tim/gits/sky130_ef_ip__ccomp3v/xschem/scomp_bias.sym
** sch_path: /home/tim/gits/sky130_ef_ip__ccomp3v/xschem/scomp_bias.sch
.subckt scomp_bias VDD VSS VBN ena3v3
*.PININFO VBN:O VDD:B VSS:B ena3v3:I
XM3 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM4 net3 net1 net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM5 VBN VBN net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=15 W=1 nf=1 m=1
XM1 VBN VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM2 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM8 net3 ena3v3 VBN VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XR2 net2 VDD VSS sky130_fd_pr__res_high_po_1p41 L=135 mult=1 m=1
.ends


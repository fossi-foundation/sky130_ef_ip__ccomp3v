magic
tech sky130A
magscale 1 2
timestamp 1747681386
<< dnwell >>
rect 4 370 8564 4032
rect 4 -3044 11126 370
<< nwell >>
rect -106 3826 8674 4142
rect -106 -2838 210 3826
rect 2532 3494 7612 3826
rect 2532 3392 4940 3494
rect 4172 3060 4940 3392
rect 4730 2314 4940 3060
rect 4778 324 4940 2314
rect 8358 546 8674 3826
rect 8358 164 11236 546
rect 10920 -2838 11236 164
rect -106 -3154 11236 -2838
<< mvnsubdiff >>
rect -39 4055 8593 4075
rect -39 4021 41 4055
rect 8328 4021 8593 4055
rect -39 4001 8593 4021
rect -39 3995 35 4001
rect -39 -3007 -19 3995
rect 15 -3007 35 3995
rect 8519 3970 8593 4001
rect 8519 356 8539 3970
rect 8573 356 8593 3970
rect 8519 323 8593 356
rect 8519 303 11163 323
rect 8519 269 8632 303
rect 11050 269 11163 303
rect 8519 249 11163 269
rect 11089 220 11163 249
rect -39 -3013 35 -3007
rect 6346 -3013 6408 -2799
rect 11089 -3007 11109 220
rect 11143 -3007 11163 220
rect 11089 -3013 11163 -3007
rect -39 -3033 11163 -3013
rect -39 -3067 41 -3033
rect 11083 -3067 11163 -3033
rect -39 -3087 11163 -3067
<< mvnsubdiffcont >>
rect 41 4021 8328 4055
rect -19 -3007 15 3995
rect 8539 356 8573 3970
rect 8632 269 11050 303
rect 11109 -3007 11143 220
rect 41 -3067 11083 -3033
<< locali >>
rect -39 4061 8594 4076
rect -39 4055 60 4061
rect 8308 4055 8594 4061
rect -39 4021 41 4055
rect 8328 4021 8594 4055
rect -39 4015 60 4021
rect 8308 4015 8594 4021
rect -39 4001 8594 4015
rect -39 3995 36 4001
rect -39 3981 -19 3995
rect 15 3981 36 3995
rect -39 -2979 -25 3981
rect 17 -2979 36 3981
rect 8519 3970 8594 4001
rect 8519 3940 8539 3970
rect 8573 3940 8594 3970
rect 8519 387 8531 3940
rect 8576 387 8594 3940
rect 9365 3549 9563 3561
rect 9365 3434 9377 3549
rect 9549 3434 9563 3549
rect 9365 3423 9563 3434
rect 9368 3031 9549 3044
rect 9368 2910 9383 3031
rect 9536 2910 9549 3031
rect 9368 2899 9549 2910
rect 10040 1368 10374 1376
rect 10040 1268 10178 1368
rect 10356 1268 10374 1368
rect 10040 1258 10374 1268
rect 8519 356 8539 387
rect 8573 356 8594 387
rect 8519 324 8594 356
rect 8519 307 11164 324
rect 8519 305 10350 307
rect 8519 303 8647 305
rect 10168 303 10350 305
rect 11031 303 11164 307
rect 8519 269 8632 303
rect 11050 269 11164 303
rect 8519 262 8647 269
rect 10168 265 10350 269
rect 11031 265 11164 269
rect 10168 262 11164 265
rect 8519 249 11164 262
rect 11089 220 11164 249
rect 11089 195 11109 220
rect 11143 195 11164 220
rect 11089 -48 11102 195
rect -39 -3007 -19 -2979
rect 15 -3007 36 -2979
rect -39 -3012 36 -3007
rect 6346 -3012 6408 -2799
rect 11088 -2983 11102 -48
rect 11146 -2983 11164 195
rect 11088 -3007 11109 -2983
rect 11143 -3007 11164 -2983
rect 11088 -3012 11164 -3007
rect -39 -3030 11164 -3012
rect -39 -3033 73 -3030
rect 11062 -3033 11164 -3030
rect -39 -3067 41 -3033
rect 11083 -3067 11164 -3033
rect -39 -3072 73 -3067
rect 11062 -3072 11164 -3067
rect -39 -3087 11164 -3072
<< viali >>
rect 60 4055 8308 4061
rect 60 4021 8308 4055
rect 60 4015 8308 4021
rect -25 -2979 -19 3981
rect -19 -2979 15 3981
rect 15 -2979 17 3981
rect 8531 387 8539 3940
rect 8539 387 8573 3940
rect 8573 387 8576 3940
rect 9377 3434 9549 3549
rect 9383 2910 9536 3031
rect 10178 1268 10356 1368
rect 8647 303 10168 305
rect 10350 303 11031 307
rect 8647 269 10168 303
rect 10350 269 11031 303
rect 8647 262 10168 269
rect 10350 265 11031 269
rect 11102 -2983 11109 195
rect 11109 -2983 11143 195
rect 11143 -2983 11146 195
rect 73 -3033 11062 -3030
rect 73 -3067 11062 -3033
rect 73 -3072 11062 -3067
<< metal1 >>
rect -39 4061 8594 4076
rect -39 4015 60 4061
rect 8308 4015 8594 4061
rect -39 4001 8594 4015
rect -39 3981 36 4001
rect -39 3834 -25 3981
rect -49 3824 -25 3834
rect 17 3834 36 3981
rect 8519 3940 8594 4001
rect 17 3824 67 3834
rect 8519 3833 8531 3940
rect -49 3087 -40 3824
rect 59 3087 67 3824
rect -49 3078 -25 3087
rect -39 -2979 -25 3078
rect 17 3078 67 3087
rect 8284 3818 8531 3833
rect 8576 3833 8594 3940
rect 9363 3922 9563 4122
rect 8576 3818 8623 3833
rect 8284 3089 8300 3818
rect 8606 3089 8623 3818
rect 9055 3402 9210 3586
rect 9436 3561 9488 3922
rect 9776 3692 10026 3704
rect 9365 3549 9563 3561
rect 9365 3434 9377 3549
rect 9549 3434 9563 3549
rect 9365 3423 9563 3434
rect 8284 3078 8531 3089
rect 17 -2979 36 3078
rect 8519 387 8531 3078
rect 8576 3078 8623 3089
rect 8576 387 8594 3078
rect 9056 1356 9210 3402
rect 9436 3044 9488 3423
rect 9776 3098 9784 3692
rect 10018 3098 10026 3692
rect 9776 3088 10026 3098
rect 9368 3031 9549 3044
rect 9368 2910 9383 3031
rect 9536 2910 9549 3031
rect 9368 2899 9549 2910
rect 9690 3012 9748 3028
rect 9436 2896 9488 2899
rect 9690 2792 9748 2806
rect 9056 1088 9212 1356
rect 9780 1350 10022 3088
rect 10160 1368 10494 1376
rect 10160 1268 10178 1368
rect 10356 1268 10494 1368
rect 10592 1358 10744 3586
rect 10160 1258 10494 1268
rect 9056 720 9062 1088
rect 9206 720 9212 1088
rect 9056 705 9212 720
rect 8519 324 8594 387
rect 8519 305 10196 324
rect 8519 262 8647 305
rect 10168 262 10196 305
rect 8519 249 10196 262
rect 10247 168 10282 1258
rect 10590 1098 10744 1358
rect 10472 1088 10744 1098
rect 10472 722 10478 1088
rect 10642 722 10744 1088
rect 10472 714 10744 722
rect 10324 307 11164 324
rect 10324 265 10350 307
rect 11031 265 11164 307
rect 10324 249 11164 265
rect 4792 134 10282 168
rect 11088 195 11164 249
rect 10736 -1268 10986 -1068
rect 10736 -1628 10986 -1428
rect -39 -3012 36 -2979
rect 6334 -3012 6420 -2822
rect 11088 -2983 11102 195
rect 11146 -2983 11164 195
rect 11088 -3012 11164 -2983
rect -39 -3030 11164 -3012
rect -39 -3072 73 -3030
rect 11062 -3072 11164 -3030
rect -39 -3087 11164 -3072
<< via1 >>
rect -40 3087 -25 3824
rect -25 3087 17 3824
rect 17 3087 59 3824
rect 8300 3089 8531 3818
rect 8531 3089 8576 3818
rect 8576 3089 8606 3818
rect 9784 3098 10018 3692
rect 9690 2806 9748 3012
rect 9062 720 9206 1088
rect 10478 722 10642 1088
<< metal2 >>
rect -49 3824 10854 3834
rect -49 3087 -40 3824
rect 59 3818 10854 3824
rect 59 3089 8300 3818
rect 8606 3692 10854 3818
rect 8606 3098 9784 3692
rect 10018 3098 10854 3692
rect 8606 3089 10854 3098
rect 59 3087 10854 3089
rect -49 3078 10854 3087
rect 8247 2806 9690 3012
rect 9748 2806 10854 3012
rect 10652 1736 10852 1792
rect 8046 1636 10852 1736
rect 10652 1592 10852 1636
rect 8288 1088 10854 1096
rect 8288 720 9062 1088
rect 9206 722 10478 1088
rect 10642 722 10854 1088
rect 9206 720 10854 722
rect 8288 714 10854 720
rect -61 -2786 6153 -2078
rect 6200 -2659 6555 -2077
rect 6199 -2787 6555 -2659
rect 6670 -2786 10764 -2658
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 1 9087 -1 0 3652
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 -1 10715 1 0 3460
box -66 -43 258 897
use comparator_high_gain  x1
timestamp 1747681386
transform -1 0 11226 0 1 438
box 69 -3444 7124 3348
use scomp_bias  x2
timestamp 1731032193
transform -1 0 5269 0 1 -1439
box 323 -1349 5039 5225
use sky130_fd_sc_hvl__lsbuflv2hv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1746753973
transform 0 1 9087 -1 0 3460
box -66 -43 2178 1671
<< labels >>
flabel metal1 10736 -1628 10936 -1428 0 FreeSans 256 0 0 0 VINM
port 6 nsew
flabel metal1 10736 -1268 10936 -1068 0 FreeSans 256 0 0 0 VINP
port 5 nsew
flabel metal2 6305 -2511 6505 -2311 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 9363 3922 9563 4122 0 FreeSans 256 0 0 0 ENA
port 7 nsew
flabel metal2 10652 1592 10852 1792 0 FreeSans 256 0 0 0 VOUT
port 0 nsew
flabel metal2 10654 808 10854 1008 0 FreeSans 256 0 0 0 DVSS
port 2 nsew
flabel metal2 10650 2806 10850 3006 0 FreeSans 256 0 0 0 DVDD
port 1 nsew
flabel metal2 10632 3516 10832 3716 0 FreeSans 256 0 0 0 VDD
port 3 nsew
<< end >>

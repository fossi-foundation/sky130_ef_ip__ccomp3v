magic
tech sky130A
magscale 1 2
timestamp 1747681611
<< dnwell >>
rect -132 -2510 11126 10125
<< nwell >>
rect -241 10017 11235 10234
rect -241 7975 76 10017
rect -241 5932 74 7975
rect 10224 6187 11235 10017
rect -241 1870 94 5932
rect 5141 5929 11235 6187
rect 9361 5860 11235 5929
rect 10900 1870 11235 5860
rect -241 -2304 74 1870
rect 10920 -2304 11235 1870
rect -241 -2619 11235 -2304
<< mvpsubdiff >>
rect -363 10323 -303 10357
rect 11302 10323 11362 10357
rect -363 10297 -329 10323
rect 11328 10297 11362 10323
rect -363 -2710 -329 -2684
rect 11328 -2710 11362 -2684
rect -363 -2744 -303 -2710
rect 11302 -2744 11362 -2710
<< mvnsubdiff >>
rect -175 10148 11169 10168
rect -175 10114 -95 10148
rect 11089 10114 11169 10148
rect -175 10094 11169 10114
rect -175 10088 -101 10094
rect -175 -2473 -155 10088
rect -121 -2473 -101 10088
rect -175 -2479 -101 -2473
rect 11095 10088 11169 10094
rect 11095 5833 11115 10088
rect 11149 5833 11169 10088
rect 11095 5785 11169 5833
rect 11095 5730 11115 5785
rect 11149 5730 11169 5785
rect 11095 5575 11169 5730
rect 11095 -2464 11115 5575
rect 11149 -2464 11169 5575
rect 11095 -2479 11169 -2464
rect -175 -2499 11169 -2479
rect -175 -2533 -95 -2499
rect 11079 -2533 11169 -2499
rect -175 -2553 11169 -2533
<< mvpsubdiffcont >>
rect -303 10323 11302 10357
rect -363 -2684 -329 10297
rect 11328 -2684 11362 10297
rect -303 -2744 11302 -2710
<< mvnsubdiffcont >>
rect -95 10114 11089 10148
rect -155 -2473 -121 10088
rect 11115 5833 11149 10088
rect 11115 5730 11149 5785
rect 11115 -2464 11149 5575
rect -95 -2533 11079 -2499
<< locali >>
rect -363 10323 -303 10357
rect 11302 10323 11362 10357
rect -363 10317 11362 10323
rect -363 10297 -221 10317
rect -329 10268 -221 10297
rect 11200 10297 11362 10317
rect 11200 10268 11328 10297
rect -329 10235 11328 10268
rect -329 10154 -242 10235
rect -329 -2544 -317 10154
rect -265 -2544 -242 10154
rect 11234 10193 11328 10235
rect -155 10114 -95 10148
rect 11089 10114 11149 10148
rect -155 10088 11149 10114
rect -121 10065 11115 10088
rect -121 10015 43 10065
rect 10930 10015 11115 10065
rect -121 9970 11115 10015
rect -121 9936 22 9970
rect -121 -2339 -100 9936
rect -46 -2339 22 9936
rect 10960 9915 11115 9970
rect 10960 5851 11005 9915
rect 11057 5851 11115 9915
rect 10960 5833 11115 5851
rect -121 -2344 22 -2339
rect 10959 5785 11149 5833
rect 10959 5730 11115 5785
rect 10959 5713 11149 5730
rect 10959 -2344 11005 5713
rect -121 -2351 11005 -2344
rect 11061 5575 11149 5713
rect 11061 -2351 11115 5575
rect -121 -2406 11115 -2351
rect -121 -2459 -9 -2406
rect 10954 -2459 11115 -2406
rect -121 -2464 11115 -2459
rect -121 -2473 11149 -2464
rect -155 -2499 11149 -2473
rect -155 -2533 -95 -2499
rect 11079 -2533 11149 -2499
rect -329 -2620 -242 -2544
rect 11234 -2592 11262 10193
rect 11319 -2592 11328 10193
rect 11234 -2620 11328 -2592
rect -329 -2649 11328 -2620
rect -329 -2684 -194 -2649
rect -363 -2689 -194 -2684
rect 11209 -2684 11328 -2649
rect 11209 -2689 11362 -2684
rect -363 -2710 11362 -2689
rect -363 -2744 -303 -2710
rect 11302 -2744 11362 -2710
<< viali >>
rect -221 10268 11200 10317
rect -317 -2544 -265 10154
rect 43 10015 10930 10065
rect -100 -2339 -46 9936
rect 11005 5851 11057 9915
rect 11005 -2351 11061 5713
rect -9 -2459 10954 -2406
rect 11262 -2592 11319 10193
rect -194 -2689 11209 -2649
<< metal1 >>
rect -363 10317 11362 10357
rect -363 10268 -221 10317
rect 11200 10268 11362 10317
rect -363 10235 11362 10268
rect -363 10154 -242 10235
rect -363 -2544 -317 10154
rect -265 -2544 -242 10154
rect 11234 10193 11362 10235
rect -113 10065 11075 10085
rect -113 10015 43 10065
rect 10930 10015 11075 10065
rect -113 10002 11075 10015
rect -113 9936 -30 10002
rect 5161 9987 5347 10002
rect -113 -2339 -100 9936
rect -46 -2339 -30 9936
rect 10992 9915 11075 10002
rect 10992 6175 11005 9915
rect 10866 6164 11005 6175
rect 11057 6175 11075 9915
rect 11234 7635 11262 10193
rect 11162 7627 11262 7635
rect 11319 7627 11362 10193
rect 11057 6164 11097 6175
rect 10866 5944 10900 6164
rect 11086 5944 11097 6164
rect 10866 5935 11005 5944
rect -113 -2388 -30 -2339
rect 10992 5851 11005 5935
rect 11057 5936 11097 5944
rect 11057 5935 11088 5936
rect 11057 5851 11075 5935
rect 11334 5899 11362 7627
rect 11162 5891 11262 5899
rect 10992 5713 11075 5851
rect 10992 -2351 11005 5713
rect 11061 -2351 11075 5713
rect 10992 -2388 11075 -2351
rect -113 -2406 11075 -2388
rect -113 -2459 -9 -2406
rect 10954 -2459 11075 -2406
rect -113 -2471 11075 -2459
rect -363 -2574 -242 -2544
rect -363 -2620 3257 -2574
rect 11234 -2592 11262 5891
rect 11319 -2592 11362 5899
rect 11234 -2620 11362 -2592
rect -363 -2649 11362 -2620
rect -363 -2689 -194 -2649
rect 11209 -2689 11362 -2649
rect -363 -2744 11362 -2689
rect -360 -2797 3257 -2744
<< via1 >>
rect 10900 5944 11005 6164
rect 11005 5944 11057 6164
rect 11057 5944 11086 6164
rect 11162 5899 11262 7627
rect 11262 5899 11319 7627
rect 11319 5899 11334 7627
<< metal2 >>
rect 5161 9987 5347 10085
rect 11138 7627 11361 7653
rect 4961 6175 5147 6257
rect 9712 6164 11097 6175
rect 9712 6163 10900 6164
rect 9712 5949 9725 6163
rect 10824 5949 10900 6163
rect 9712 5944 10900 5949
rect 11086 5944 11097 6164
rect 9712 5936 11097 5944
rect 9712 5935 11088 5936
rect 4961 5914 5147 5935
rect 11138 5899 11162 7627
rect 11334 5899 11361 7627
rect 11138 4077 11361 5899
rect 10640 3417 11362 3922
rect -181 1871 198 1971
rect 10922 1738 11362 1838
rect -181 1636 198 1736
<< via2 >>
rect 4961 5935 5147 6175
rect 9725 5949 10824 6163
<< metal3 >>
rect 623 2142 723 7084
rect 1659 6114 1759 7545
rect 4954 6175 5158 6184
rect 835 6014 1759 6114
rect 2077 6160 4961 6175
rect 835 1343 935 6014
rect 2077 5948 2090 6160
rect 2488 5948 4961 6160
rect 2077 5935 4961 5948
rect 5147 6163 11039 6175
rect 5147 5949 9725 6163
rect 10824 5949 11039 6163
rect 5147 5935 11039 5949
rect 4954 5927 5158 5935
<< via3 >>
rect 2090 5948 2488 6160
<< metal4 >>
rect 285 9775 1485 10036
rect 2570 9770 3770 10036
rect 285 6171 1485 6273
rect 2769 6216 6781 6936
rect 1685 6171 2501 6173
rect 285 6160 2501 6171
rect 285 5948 2090 6160
rect 2488 5948 2501 6160
rect 285 4660 2501 5948
rect 6061 5601 6781 6216
use cc_via2_3cut  cc_via2_3cut_0
timestamp 1717772055
transform 0 1 -639040 -1 0 518654
box 517199 639873 517310 640172
use cc_via2_3cut  cc_via2_3cut_1
timestamp 1717772055
transform 0 1 -639448 -1 0 519454
box 517199 639873 517310 640172
use comparator_bias  comparator_bias_0
timestamp 1747681611
transform -1 0 518254 0 1 -639855
box 508008 646042 518182 649916
use comparator_core  comparator_core_0
timestamp 1718227246
transform 1 0 -506140 0 1 -641069
box 506214 638825 517124 647001
<< labels >>
flabel metal2 -140 1636 198 1736 0 FreeSans 1600 0 0 0 VINM
port 0 nsew
flabel metal2 -140 1871 198 1971 0 FreeSans 1600 0 0 0 VINP
port 1 nsew
flabel metal4 2570 9770 3770 10036 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
flabel metal4 285 9775 1485 10036 0 FreeSans 1600 0 0 0 VDD
port 2 nsew
flabel metal2 10927 3417 11362 3922 0 FreeSans 1600 0 0 0 DVDD
port 5 nsew
flabel metal2 10936 1738 11362 1838 0 FreeSans 1200 0 0 0 VOUT
port 7 nsew
flabel metal2 11138 4077 11361 5865 0 FreeSans 1600 270 0 0 DVSS
port 6 nsew
<< end >>
